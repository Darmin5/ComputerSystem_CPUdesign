module count10_tb(

    );
    reg rst;
    reg clk;
    reg en;
    wire [3:0] count;
    wire co;
    initial begin
        rst = 0;
        clk = 0;
        en = 0;
        #10
        rst = 1;
        #10
        rst = 0;
        en = 1;
    end
    
    always #10 clk = ~clk;
    count_10 count10(rst,clk,en,count,co);    
endmodule
